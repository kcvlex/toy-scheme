`default_nettype none

module top();
    reg CLK, RST_X;
    initial begin CLK = 1; forever #50 CLK = ~CLK; end
    initial begin RST_X = 0; #125 RST_X = 1;       end
    initial begin p.PC = 4; end
    initial begin #10000 $finish(); end
    initial begin $dumpfile("wave.vcd"); $dumpvars(0, p); end

    initial begin
        /*
        p.imem.mem[0] = 32'd0;
        p.imem.mem[1] = { 12'd10, 5'd0, 3'b0, 5'd5, 7'b0010011 };
        p.imem.mem[2] = { 12'd32, 5'd0, 3'b0, 5'd6, 7'b0010011 };
        p.imem.mem[3] = { 7'd0, 5'd6, 5'd5, 3'b0, 5'd7, 7'b0110011 };
        */

        /*
        // -42 + 48
        p.imem.mem[0] = 32'd0;
        p.imem.mem[1] = 32'b11111101000000000000001010010011;
        p.imem.mem[2] = 32'b00000010101000000000001100010011;
        p.imem.mem[3] = 32'b00000000011000101000001110110011;
        */
p.imem.mem[0] = 32'b00000000000000000000000000010011;
p.imem.mem[1] = 32'b00000000000000000000000000010011;
p.imem.mem[2] = 32'b00000000000000000000000000010011;
p.imem.mem[3] = 32'b00001110100000000000000011101111;
p.imem.mem[4] = 32'b00000000000000000110000010110011;
p.imem.mem[5] = 32'b00000000000000001000000001100111;
p.imem.mem[6] = 32'b00000000001000010010000000100011;
p.imem.mem[7] = 32'b11111111110000010000000100010011;
p.imem.mem[8] = 32'b00000000000100010010000000100011;
p.imem.mem[9] = 32'b11111111110000010000000100010011;
p.imem.mem[10] = 32'b00000000100000010010000000100011;
p.imem.mem[11] = 32'b11111111110000010000000100010011;
p.imem.mem[12] = 32'b00000000001000010110010000110011;
p.imem.mem[13] = 32'b00000000101000010010000000100011;
p.imem.mem[14] = 32'b11111111110000010000000100010011;
p.imem.mem[15] = 32'b00000000110001100110010100110011;
p.imem.mem[16] = 32'b00000000101000010010000000100011;
p.imem.mem[17] = 32'b11111111110000010000000100010011;
p.imem.mem[18] = 32'b00000000101000010010000000100011;
p.imem.mem[19] = 32'b11111111110000010000000100010011;
p.imem.mem[20] = 32'b00000000110101101110010100110011;
p.imem.mem[21] = 32'b00000000101000010010000000100011;
p.imem.mem[22] = 32'b11111111110000010000000100010011;
p.imem.mem[23] = 32'b00000000101000010010000000100011;
p.imem.mem[24] = 32'b11111111110000010000000100010011;
p.imem.mem[25] = 32'b00000000000100000000010100010011;
p.imem.mem[26] = 32'b00000000101000010010000000100011;
p.imem.mem[27] = 32'b11111111110000010000000100010011;
p.imem.mem[28] = 32'b00000000001000000000010100010011;
p.imem.mem[29] = 32'b00000000101000010010000000100011;
p.imem.mem[30] = 32'b11111111110000010000000100010011;
p.imem.mem[31] = 32'b00000000010000010010001110000011;
p.imem.mem[32] = 32'b00000000010000010000000100010011;
p.imem.mem[33] = 32'b00000000010000010010001100000011;
p.imem.mem[34] = 32'b00000000010000010000000100010011;
p.imem.mem[35] = 32'b00000000010000010010010100000011;
p.imem.mem[36] = 32'b00000000010000010000000100010011;
p.imem.mem[37] = 32'b00000000011100110000010100110011;
p.imem.mem[38] = 32'b00000000101000010010000000100011;
p.imem.mem[39] = 32'b11111111110000010000000100010011;
p.imem.mem[40] = 32'b00000000010000010010001110000011;
p.imem.mem[41] = 32'b00000000010000010000000100010011;
p.imem.mem[42] = 32'b00000000010000010010001100000011;
p.imem.mem[43] = 32'b00000000010000010000000100010011;
p.imem.mem[44] = 32'b00000000010000010010010100000011;
p.imem.mem[45] = 32'b00000000010000010000000100010011;
p.imem.mem[46] = 32'b00000000011100110000010100110011;
p.imem.mem[47] = 32'b00000000101000010010000000100011;
p.imem.mem[48] = 32'b11111111110000010000000100010011;
p.imem.mem[49] = 32'b00000000010000010010001110000011;
p.imem.mem[50] = 32'b00000000010000010000000100010011;
p.imem.mem[51] = 32'b00000000010000010010001100000011;
p.imem.mem[52] = 32'b00000000010000010000000100010011;
p.imem.mem[53] = 32'b00000000010000010010010100000011;
p.imem.mem[54] = 32'b00000000010000010000000100010011;
p.imem.mem[55] = 32'b00000000011100110000010100110011;
p.imem.mem[56] = 32'b00000000100001000110001010110011;
p.imem.mem[57] = 32'b00000000110000101010000010000011;
p.imem.mem[58] = 32'b00000000100000101010000100000011;
p.imem.mem[59] = 32'b00000000010000101010010000000011;
p.imem.mem[60] = 32'b00000000000000001000000001100111;
p.imem.mem[61] = 32'b00000000101000010010000000100011;
p.imem.mem[62] = 32'b11111111110000010000000100010011;
p.imem.mem[63] = 32'b00000000000100010010000000100011;
p.imem.mem[64] = 32'b11111111110000010000000100010011;
p.imem.mem[65] = 32'b00000010110000000000010100010011;
p.imem.mem[66] = 32'b00000000101001010110011010110011;
p.imem.mem[67] = 32'b00000010101100000000010100010011;
p.imem.mem[68] = 32'b00000000101001010110011000110011;
p.imem.mem[69] = 32'b00000010101000000000010100010011;
p.imem.mem[70] = 32'b00000000101001010110010110110011;
p.imem.mem[71] = 32'b00000000010000010010000000000011;
p.imem.mem[72] = 32'b00000000010000010000000100010011;
p.imem.mem[73] = 32'b11101111010111111111000011101111;
p.imem.mem[74] = 32'b00000000010000010010000010000011;
p.imem.mem[75] = 32'b00000000010000010000000100010011;
end
always @(p.PC) begin if (p.PC[11:2] == 0) $finish(); end
    
    always @(CLK) begin
        #30 $write("%d : %d \t %d %d %d %d \t %d %d %d %b \t %d %d %d \t %d %d %d %d %d \t %b\n",
                $stime-30, 
                p.PC,
                p.cpu.rs1, p.cpu.rs2, p.cpu.rd, $signed(p.cpu.imm),
                $signed(p.cpu.rrs1), $signed(p.cpu.rrs2), $signed(p.cpu.Ex_wd_mem), $signed(p.cpu.Ex_store),
                $signed(p.cpu.alu_cont.alu.lhs), $signed(p.cpu.alu_cont.alu.rhs), $signed(p.cpu.alu_cont.alu.res),
                $signed(p.cpu.regfile.x[6]), $signed(p.cpu.regfile.x[7]), $signed(p.cpu.regfile.x[10]), $signed(p.cpu.regfile.x[11]), $signed(p.cpu.regfile.x[1]),
                p.cpu.instr_type);
    end

    PROCESSOR p(CLK, RST_X);
endmodule


module PROCESSOR(
    input wire CLK,
    input wire RST_X
);
    reg [31:0] PC;
    wire [31:0] instr, next_pc;

    always @(posedge RST_X) PC <= #1 4;
    always @(posedge CLK) if (RST_X) PC <= #1 next_pc;

    IMEM imem(CLK, RST_X, PC, instr);
    CPU cpu(CLK, RST_X, PC, instr, next_pc);
endmodule
